library verilog;
use verilog.vl_types.all;
entity Interface is
end Interface;
